library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity tuberom_65c102 is
    port (
        CLK  : in  std_logic;
        ADDR : in  std_logic_vector(10 downto 0);
        DATA : out std_logic_vector(7 downto 0)
        );
end;

architecture RTL of tuberom_65c102 is

    type rom_t is array(0 to  2047) of std_logic_vector(7 downto 0);
    signal rom : rom_t := (
             x"A2",
             x"00",
             x"BD",
             x"00",
             x"FF",
             x"9D",
             x"00",
             x"FF",
             x"CA",
             x"D0",
             x"F7",
             x"A2",
             x"36",
             x"BD",
             x"80",
             x"FF",
             x"9D",
             x"00",
             x"02",
             x"CA",
             x"10",
             x"F7",
             x"9A",
             x"A2",
             x"F0",
             x"BD",
             x"FF",
             x"FD",
             x"9D",
             x"FF",
             x"FD",
             x"CA",
             x"D0",
             x"F7",
             x"A0",
             x"00",
             x"84",
             x"F8",
             x"A9",
             x"F8",
             x"85",
             x"F9",
             x"B1",
             x"F8",
             x"91",
             x"F8",
             x"C8",
             x"D0",
             x"F9",
             x"E6",
             x"F9",
             x"A5",
             x"F9",
             x"C9",
             x"FE",
             x"D0",
             x"F1",
             x"A2",
             x"10",
             x"BD",
             x"59",
             x"F8",
             x"9D",
             x"00",
             x"01",
             x"CA",
             x"10",
             x"F7",
             x"A5",
             x"EE",
             x"85",
             x"F6",
             x"A5",
             x"EF",
             x"85",
             x"F7",
             x"A9",
             x"00",
             x"85",
             x"FF",
             x"85",
             x"F2",
             x"A9",
             x"F8",
             x"85",
             x"F3",
             x"4C",
             x"00",
             x"01",
             x"AD",
             x"F8",
             x"FE",
             x"58",
             x"4C",
             x"60",
             x"F8",
             x"20",
             x"A5",
             x"FE",
             x"0A",
             x"41",
             x"63",
             x"6F",
             x"72",
             x"6E",
             x"20",
             x"54",
             x"55",
             x"42",
             x"45",
             x"20",
             x"36",
             x"35",
             x"43",
             x"31",
             x"30",
             x"32",
             x"20",
             x"43",
             x"6F",
             x"2D",
             x"50",
             x"72",
             x"6F",
             x"63",
             x"65",
             x"73",
             x"73",
             x"6F",
             x"72",
             x"0A",
             x"0A",
             x"0D",
             x"00",
             x"EA",
             x"A9",
             x"98",
             x"8D",
             x"5E",
             x"F8",
             x"A9",
             x"F8",
             x"8D",
             x"5F",
             x"F8",
             x"20",
             x"80",
             x"F9",
             x"C9",
             x"80",
             x"F0",
             x"28",
             x"A9",
             x"2A",
             x"20",
             x"EE",
             x"FF",
             x"A2",
             x"68",
             x"A0",
             x"F9",
             x"A9",
             x"00",
             x"20",
             x"F1",
             x"FF",
             x"B0",
             x"0A",
             x"A2",
             x"36",
             x"A0",
             x"02",
             x"20",
             x"F7",
             x"FF",
             x"4C",
             x"98",
             x"F8",
             x"A9",
             x"7E",
             x"20",
             x"F4",
             x"FF",
             x"00",
             x"11",
             x"45",
             x"73",
             x"63",
             x"61",
             x"70",
             x"65",
             x"00",
             x"A5",
             x"F6",
             x"85",
             x"EE",
             x"85",
             x"F2",
             x"A5",
             x"F7",
             x"85",
             x"EF",
             x"85",
             x"F3",
             x"A0",
             x"07",
             x"B1",
             x"EE",
             x"D8",
             x"18",
             x"65",
             x"EE",
             x"85",
             x"FD",
             x"A9",
             x"00",
             x"65",
             x"EF",
             x"85",
             x"FE",
             x"A0",
             x"00",
             x"B1",
             x"FD",
             x"D0",
             x"23",
             x"C8",
             x"B1",
             x"FD",
             x"C9",
             x"28",
             x"D0",
             x"1C",
             x"C8",
             x"B1",
             x"FD",
             x"C9",
             x"43",
             x"D0",
             x"15",
             x"C8",
             x"B1",
             x"FD",
             x"C9",
             x"29",
             x"D0",
             x"0E",
             x"A0",
             x"06",
             x"B1",
             x"EE",
             x"29",
             x"4F",
             x"C9",
             x"40",
             x"90",
             x"09",
             x"29",
             x"0D",
             x"D0",
             x"28",
             x"A9",
             x"01",
             x"6C",
             x"F2",
             x"00",
             x"A9",
             x"50",
             x"8D",
             x"02",
             x"02",
             x"A9",
             x"F9",
             x"8D",
             x"03",
             x"02",
             x"00",
             x"00",
             x"54",
             x"68",
             x"69",
             x"73",
             x"20",
             x"69",
             x"73",
             x"20",
             x"6E",
             x"6F",
             x"74",
             x"20",
             x"61",
             x"20",
             x"6C",
             x"61",
             x"6E",
             x"67",
             x"75",
             x"61",
             x"67",
             x"65",
             x"00",
             x"A9",
             x"50",
             x"8D",
             x"02",
             x"02",
             x"A9",
             x"F9",
             x"8D",
             x"03",
             x"02",
             x"00",
             x"00",
             x"49",
             x"20",
             x"63",
             x"61",
             x"6E",
             x"6E",
             x"6F",
             x"74",
             x"20",
             x"72",
             x"75",
             x"6E",
             x"20",
             x"74",
             x"68",
             x"69",
             x"73",
             x"20",
             x"63",
             x"6F",
             x"64",
             x"65",
             x"00",
             x"A2",
             x"FF",
             x"9A",
             x"20",
             x"E7",
             x"FF",
             x"A0",
             x"01",
             x"B1",
             x"FD",
             x"F0",
             x"06",
             x"20",
             x"EE",
             x"FF",
             x"C8",
             x"D0",
             x"F6",
             x"20",
             x"E7",
             x"FF",
             x"4C",
             x"98",
             x"F8",
             x"36",
             x"02",
             x"CA",
             x"20",
             x"FF",
             x"2C",
             x"F8",
             x"FE",
             x"EA",
             x"50",
             x"FA",
             x"8D",
             x"F9",
             x"FE",
             x"60",
             x"A9",
             x"00",
             x"20",
             x"57",
             x"FC",
             x"20",
             x"80",
             x"F9",
             x"0A",
             x"2C",
             x"FA",
             x"FE",
             x"10",
             x"FB",
             x"AD",
             x"FB",
             x"FE",
             x"60",
             x"C8",
             x"B1",
             x"F8",
             x"C9",
             x"20",
             x"F0",
             x"F9",
             x"60",
             x"A2",
             x"00",
             x"86",
             x"F0",
             x"86",
             x"F1",
             x"B1",
             x"F8",
             x"C9",
             x"30",
             x"90",
             x"1F",
             x"C9",
             x"3A",
             x"90",
             x"0A",
             x"29",
             x"DF",
             x"E9",
             x"07",
             x"90",
             x"15",
             x"C9",
             x"40",
             x"B0",
             x"11",
             x"0A",
             x"0A",
             x"0A",
             x"0A",
             x"A2",
             x"03",
             x"0A",
             x"26",
             x"F0",
             x"26",
             x"F1",
             x"CA",
             x"10",
             x"F8",
             x"C8",
             x"D0",
             x"DB",
             x"60",
             x"86",
             x"F8",
             x"84",
             x"F9",
             x"A0",
             x"00",
             x"2C",
             x"FA",
             x"FE",
             x"50",
             x"FB",
             x"B1",
             x"F8",
             x"8D",
             x"FB",
             x"FE",
             x"C8",
             x"C9",
             x"0D",
             x"D0",
             x"F1",
             x"A4",
             x"F9",
             x"60",
             x"48",
             x"86",
             x"F8",
             x"84",
             x"F9",
             x"A0",
             x"00",
             x"20",
             x"8A",
             x"F9",
             x"C8",
             x"C9",
             x"2A",
             x"F0",
             x"F8",
             x"29",
             x"DF",
             x"AA",
             x"B1",
             x"F8",
             x"E0",
             x"47",
             x"F0",
             x"5E",
             x"E0",
             x"48",
             x"D0",
             x"49",
             x"C9",
             x"2E",
             x"F0",
             x"2D",
             x"29",
             x"DF",
             x"C9",
             x"45",
             x"D0",
             x"3F",
             x"C8",
             x"B1",
             x"F8",
             x"C9",
             x"2E",
             x"F0",
             x"20",
             x"29",
             x"DF",
             x"C9",
             x"4C",
             x"D0",
             x"32",
             x"C8",
             x"B1",
             x"F8",
             x"C9",
             x"2E",
             x"F0",
             x"13",
             x"29",
             x"DF",
             x"C9",
             x"50",
             x"D0",
             x"25",
             x"C8",
             x"B1",
             x"F8",
             x"29",
             x"DF",
             x"C9",
             x"41",
             x"90",
             x"04",
             x"C9",
             x"5B",
             x"90",
             x"18",
             x"20",
             x"A5",
             x"FE",
             x"0A",
             x"0D",
             x"36",
             x"35",
             x"43",
             x"31",
             x"30",
             x"32",
             x"20",
             x"54",
             x"55",
             x"42",
             x"45",
             x"20",
             x"31",
             x"2E",
             x"31",
             x"30",
             x"0A",
             x"0D",
             x"EA",
             x"A9",
             x"02",
             x"20",
             x"57",
             x"FC",
             x"20",
             x"C1",
             x"F9",
             x"20",
             x"80",
             x"F9",
             x"C9",
             x"80",
             x"F0",
             x"20",
             x"68",
             x"60",
             x"29",
             x"DF",
             x"C9",
             x"4F",
             x"D0",
             x"E9",
             x"20",
             x"89",
             x"F9",
             x"20",
             x"91",
             x"F9",
             x"20",
             x"8A",
             x"F9",
             x"C9",
             x"0D",
             x"D0",
             x"DC",
             x"8A",
             x"F0",
             x"08",
             x"A5",
             x"F0",
             x"85",
             x"F6",
             x"A5",
             x"F1",
             x"85",
             x"F7",
             x"A5",
             x"EF",
             x"48",
             x"A5",
             x"EE",
             x"48",
             x"20",
             x"C0",
             x"F8",
             x"68",
             x"85",
             x"EE",
             x"85",
             x"F2",
             x"68",
             x"85",
             x"EF",
             x"85",
             x"F3",
             x"68",
             x"60",
             x"F0",
             x"C2",
             x"C9",
             x"80",
             x"B0",
             x"25",
             x"48",
             x"A9",
             x"04",
             x"2C",
             x"FA",
             x"FE",
             x"50",
             x"FB",
             x"8D",
             x"FB",
             x"FE",
             x"2C",
             x"FA",
             x"FE",
             x"50",
             x"FB",
             x"8E",
             x"FB",
             x"FE",
             x"68",
             x"2C",
             x"FA",
             x"FE",
             x"50",
             x"FB",
             x"8D",
             x"FB",
             x"FE",
             x"2C",
             x"FA",
             x"FE",
             x"10",
             x"FB",
             x"AE",
             x"FB",
             x"FE",
             x"60",
             x"C9",
             x"82",
             x"F0",
             x"5A",
             x"C9",
             x"83",
             x"F0",
             x"51",
             x"C9",
             x"84",
             x"F0",
             x"48",
             x"48",
             x"A9",
             x"06",
             x"2C",
             x"FA",
             x"FE",
             x"50",
             x"FB",
             x"8D",
             x"FB",
             x"FE",
             x"2C",
             x"FA",
             x"FE",
             x"50",
             x"FB",
             x"8E",
             x"FB",
             x"FE",
             x"2C",
             x"FA",
             x"FE",
             x"50",
             x"FB",
             x"8C",
             x"FB",
             x"FE",
             x"68",
             x"2C",
             x"FA",
             x"FE",
             x"50",
             x"FB",
             x"8D",
             x"FB",
             x"FE",
             x"C9",
             x"8E",
             x"F0",
             x"A1",
             x"C9",
             x"9D",
             x"F0",
             x"1B",
             x"48",
             x"2C",
             x"FA",
             x"FE",
             x"10",
             x"FB",
             x"AD",
             x"FB",
             x"FE",
             x"0A",
             x"68",
             x"2C",
             x"FA",
             x"FE",
             x"10",
             x"FB",
             x"AC",
             x"FB",
             x"FE",
             x"2C",
             x"FA",
             x"FE",
             x"10",
             x"FB",
             x"AE",
             x"FB",
             x"FE",
             x"60",
             x"A6",
             x"F2",
             x"A4",
             x"F3",
             x"60",
             x"A2",
             x"00",
             x"A0",
             x"08",
             x"60",
             x"A2",
             x"00",
             x"A0",
             x"00",
             x"60",
             x"86",
             x"F8",
             x"84",
             x"F9",
             x"A8",
             x"F0",
             x"71",
             x"48",
             x"A0",
             x"08",
             x"2C",
             x"FA",
             x"FE",
             x"50",
             x"FB",
             x"8C",
             x"FB",
             x"FE",
             x"2C",
             x"FA",
             x"FE",
             x"50",
             x"FB",
             x"8D",
             x"FB",
             x"FE",
             x"AA",
             x"10",
             x"08",
             x"A0",
             x"00",
             x"B1",
             x"F8",
             x"A8",
             x"4C",
             x"3A",
             x"FB",
             x"BC",
             x"C9",
             x"FC",
             x"E0",
             x"15",
             x"90",
             x"02",
             x"A0",
             x"10",
             x"2C",
             x"FA",
             x"FE",
             x"50",
             x"FB",
             x"8C",
             x"FB",
             x"FE",
             x"88",
             x"30",
             x"0D",
             x"2C",
             x"FA",
             x"FE",
             x"50",
             x"FB",
             x"B1",
             x"F8",
             x"8D",
             x"FB",
             x"FE",
             x"88",
             x"10",
             x"F3",
             x"8A",
             x"10",
             x"08",
             x"A0",
             x"01",
             x"B1",
             x"F8",
             x"A8",
             x"4C",
             x"66",
             x"FB",
             x"BC",
             x"DD",
             x"FC",
             x"E0",
             x"15",
             x"90",
             x"02",
             x"A0",
             x"10",
             x"2C",
             x"FA",
             x"FE",
             x"50",
             x"FB",
             x"8C",
             x"FB",
             x"FE",
             x"88",
             x"30",
             x"0D",
             x"2C",
             x"FA",
             x"FE",
             x"10",
             x"FB",
             x"AD",
             x"FB",
             x"FE",
             x"91",
             x"F8",
             x"88",
             x"10",
             x"F3",
             x"A4",
             x"F9",
             x"A6",
             x"F8",
             x"68",
             x"60",
             x"A9",
             x"0A",
             x"20",
             x"57",
             x"FC",
             x"A0",
             x"04",
             x"2C",
             x"FA",
             x"FE",
             x"50",
             x"FB",
             x"B1",
             x"F8",
             x"8D",
             x"FB",
             x"FE",
             x"88",
             x"C0",
             x"01",
             x"D0",
             x"F1",
             x"A9",
             x"07",
             x"20",
             x"57",
             x"FC",
             x"B1",
             x"F8",
             x"48",
             x"88",
             x"2C",
             x"FA",
             x"FE",
             x"50",
             x"FB",
             x"8C",
             x"FB",
             x"FE",
             x"B1",
             x"F8",
             x"48",
             x"A2",
             x"FF",
             x"20",
             x"80",
             x"F9",
             x"C9",
             x"80",
             x"B0",
             x"1D",
             x"68",
             x"85",
             x"F8",
             x"68",
             x"85",
             x"F9",
             x"A0",
             x"00",
             x"2C",
             x"FA",
             x"FE",
             x"10",
             x"FB",
             x"AD",
             x"FB",
             x"FE",
             x"91",
             x"F8",
             x"C8",
             x"C9",
             x"0D",
             x"D0",
             x"F1",
             x"A9",
             x"00",
             x"88",
             x"18",
             x"E8",
             x"60",
             x"68",
             x"68",
             x"A9",
             x"00",
             x"60",
             x"48",
             x"A9",
             x"0C",
             x"20",
             x"57",
             x"FC",
             x"2C",
             x"FA",
             x"FE",
             x"50",
             x"FB",
             x"8C",
             x"FB",
             x"FE",
             x"B5",
             x"03",
             x"20",
             x"57",
             x"FC",
             x"B5",
             x"02",
             x"20",
             x"57",
             x"FC",
             x"B5",
             x"01",
             x"20",
             x"57",
             x"FC",
             x"B5",
             x"00",
             x"20",
             x"57",
             x"FC",
             x"68",
             x"20",
             x"57",
             x"FC",
             x"20",
             x"80",
             x"F9",
             x"48",
             x"20",
             x"80",
             x"F9",
             x"95",
             x"03",
             x"20",
             x"80",
             x"F9",
             x"95",
             x"02",
             x"20",
             x"80",
             x"F9",
             x"95",
             x"01",
             x"20",
             x"80",
             x"F9",
             x"95",
             x"00",
             x"68",
             x"60",
             x"48",
             x"A9",
             x"12",
             x"20",
             x"57",
             x"FC",
             x"68",
             x"20",
             x"57",
             x"FC",
             x"C9",
             x"00",
             x"D0",
             x"0A",
             x"48",
             x"98",
             x"20",
             x"57",
             x"FC",
             x"20",
             x"80",
             x"F9",
             x"68",
             x"60",
             x"20",
             x"BD",
             x"F9",
             x"4C",
             x"80",
             x"F9",
             x"A9",
             x"0E",
             x"20",
             x"57",
             x"FC",
             x"98",
             x"20",
             x"57",
             x"FC",
             x"4C",
             x"7C",
             x"F9",
             x"48",
             x"A9",
             x"10",
             x"20",
             x"57",
             x"FC",
             x"98",
             x"20",
             x"57",
             x"FC",
             x"68",
             x"20",
             x"57",
             x"FC",
             x"48",
             x"20",
             x"80",
             x"F9",
             x"68",
             x"60",
             x"2C",
             x"FA",
             x"FE",
             x"50",
             x"FB",
             x"8D",
             x"FB",
             x"FE",
             x"60",
             x"84",
             x"FB",
             x"86",
             x"FA",
             x"48",
             x"A9",
             x"14",
             x"20",
             x"57",
             x"FC",
             x"A0",
             x"11",
             x"B1",
             x"FA",
             x"20",
             x"57",
             x"FC",
             x"88",
             x"C0",
             x"01",
             x"D0",
             x"F6",
             x"88",
             x"B1",
             x"FA",
             x"AA",
             x"C8",
             x"B1",
             x"FA",
             x"A8",
             x"20",
             x"BD",
             x"F9",
             x"68",
             x"20",
             x"57",
             x"FC",
             x"20",
             x"80",
             x"F9",
             x"48",
             x"A0",
             x"11",
             x"20",
             x"80",
             x"F9",
             x"91",
             x"FA",
             x"88",
             x"C0",
             x"01",
             x"D0",
             x"F6",
             x"A4",
             x"FB",
             x"A6",
             x"FA",
             x"68",
             x"60",
             x"84",
             x"FB",
             x"86",
             x"FA",
             x"48",
             x"A9",
             x"16",
             x"20",
             x"57",
             x"FC",
             x"A0",
             x"0C",
             x"B1",
             x"FA",
             x"20",
             x"57",
             x"FC",
             x"88",
             x"10",
             x"F8",
             x"68",
             x"20",
             x"57",
             x"FC",
             x"A0",
             x"0C",
             x"20",
             x"80",
             x"F9",
             x"91",
             x"FA",
             x"88",
             x"10",
             x"F8",
             x"A4",
             x"FB",
             x"A6",
             x"FA",
             x"4C",
             x"7C",
             x"F9",
             x"00",
             x"FF",
             x"42",
             x"61",
             x"64",
             x"00",
             x"00",
             x"05",
             x"00",
             x"05",
             x"04",
             x"05",
             x"08",
             x"0E",
             x"04",
             x"01",
             x"01",
             x"05",
             x"00",
             x"01",
             x"20",
             x"10",
             x"0D",
             x"00",
             x"04",
             x"80",
             x"05",
             x"00",
             x"05",
             x"00",
             x"05",
             x"00",
             x"00",
             x"00",
             x"05",
             x"09",
             x"05",
             x"00",
             x"08",
             x"18",
             x"00",
             x"01",
             x"0D",
             x"80",
             x"04",
             x"80",
             x"85",
             x"FC",
             x"68",
             x"48",
             x"29",
             x"10",
             x"D0",
             x"10",
             x"6C",
             x"04",
             x"02",
             x"2C",
             x"FE",
             x"FE",
             x"30",
             x"4A",
             x"2C",
             x"F8",
             x"FE",
             x"30",
             x"1E",
             x"6C",
             x"06",
             x"02",
             x"8A",
             x"48",
             x"BA",
             x"BD",
             x"03",
             x"01",
             x"D8",
             x"38",
             x"E9",
             x"01",
             x"85",
             x"FD",
             x"BD",
             x"04",
             x"01",
             x"E9",
             x"00",
             x"85",
             x"FE",
             x"68",
             x"AA",
             x"A5",
             x"FC",
             x"58",
             x"6C",
             x"02",
             x"02",
             x"AD",
             x"F9",
             x"FE",
             x"30",
             x"1C",
             x"98",
             x"48",
             x"8A",
             x"48",
             x"20",
             x"8D",
             x"FE",
             x"A8",
             x"20",
             x"8D",
             x"FE",
             x"AA",
             x"20",
             x"8D",
             x"FE",
             x"20",
             x"43",
             x"FD",
             x"68",
             x"AA",
             x"68",
             x"A8",
             x"A5",
             x"FC",
             x"40",
             x"6C",
             x"20",
             x"02",
             x"0A",
             x"85",
             x"FF",
             x"A5",
             x"FC",
             x"40",
             x"AD",
             x"FF",
             x"FE",
             x"10",
             x"21",
             x"58",
             x"2C",
             x"FA",
             x"FE",
             x"10",
             x"FB",
             x"AD",
             x"FB",
             x"FE",
             x"A9",
             x"00",
             x"8D",
             x"36",
             x"02",
             x"A8",
             x"20",
             x"80",
             x"F9",
             x"8D",
             x"37",
             x"02",
             x"C8",
             x"20",
             x"80",
             x"F9",
             x"99",
             x"37",
             x"02",
             x"D0",
             x"F7",
             x"4C",
             x"36",
             x"02",
             x"8D",
             x"FA",
             x"FF",
             x"98",
             x"48",
             x"AC",
             x"FA",
             x"FF",
             x"B9",
             x"7D",
             x"FE",
             x"8D",
             x"FA",
             x"FF",
             x"B9",
             x"85",
             x"FE",
             x"8D",
             x"FB",
             x"FF",
             x"B9",
             x"6D",
             x"FE",
             x"85",
             x"F4",
             x"B9",
             x"75",
             x"FE",
             x"85",
             x"F5",
             x"2C",
             x"FE",
             x"FE",
             x"10",
             x"FB",
             x"AD",
             x"FF",
             x"FE",
             x"C0",
             x"05",
             x"F0",
             x"58",
             x"98",
             x"48",
             x"A0",
             x"01",
             x"2C",
             x"FE",
             x"FE",
             x"10",
             x"FB",
             x"AD",
             x"FF",
             x"FE",
             x"2C",
             x"FE",
             x"FE",
             x"10",
             x"FB",
             x"AD",
             x"FF",
             x"FE",
             x"2C",
             x"FE",
             x"FE",
             x"10",
             x"FB",
             x"AD",
             x"FF",
             x"FE",
             x"91",
             x"F4",
             x"88",
             x"2C",
             x"FE",
             x"FE",
             x"10",
             x"FB",
             x"AD",
             x"FF",
             x"FE",
             x"91",
             x"F4",
             x"2C",
             x"FD",
             x"FE",
             x"2C",
             x"FD",
             x"FE",
             x"2C",
             x"FE",
             x"FE",
             x"10",
             x"FB",
             x"AD",
             x"FF",
             x"FE",
             x"68",
             x"C9",
             x"06",
             x"90",
             x"1C",
             x"D0",
             x"1F",
             x"A0",
             x"00",
             x"AD",
             x"FC",
             x"FE",
             x"29",
             x"80",
             x"10",
             x"F9",
             x"B9",
             x"FF",
             x"FF",
             x"8D",
             x"FD",
             x"FE",
             x"C8",
             x"D0",
             x"F0",
             x"2C",
             x"FC",
             x"FE",
             x"10",
             x"FB",
             x"8D",
             x"FD",
             x"FE",
             x"68",
             x"A8",
             x"A5",
             x"FC",
             x"40",
             x"A0",
             x"00",
             x"AD",
             x"FC",
             x"FE",
             x"29",
             x"80",
             x"10",
             x"F9",
             x"AD",
             x"FD",
             x"FE",
             x"99",
             x"FF",
             x"FF",
             x"C8",
             x"D0",
             x"F0",
             x"F0",
             x"E7",
             x"48",
             x"AD",
             x"FF",
             x"FF",
             x"8D",
             x"FD",
             x"FE",
             x"EE",
             x"0F",
             x"FE",
             x"D0",
             x"03",
             x"EE",
             x"10",
             x"FE",
             x"68",
             x"40",
             x"48",
             x"AD",
             x"FD",
             x"FE",
             x"8D",
             x"FF",
             x"FF",
             x"EE",
             x"23",
             x"FE",
             x"D0",
             x"03",
             x"EE",
             x"24",
             x"FE",
             x"68",
             x"40",
             x"48",
             x"98",
             x"48",
             x"A0",
             x"00",
             x"B1",
             x"F6",
             x"8D",
             x"FD",
             x"FE",
             x"E6",
             x"F6",
             x"D0",
             x"02",
             x"E6",
             x"F7",
             x"B1",
             x"F6",
             x"8D",
             x"FD",
             x"FE",
             x"E6",
             x"F6",
             x"D0",
             x"02",
             x"E6",
             x"F7",
             x"68",
             x"A8",
             x"68",
             x"40",
             x"48",
             x"98",
             x"48",
             x"A0",
             x"00",
             x"AD",
             x"FD",
             x"FE",
             x"91",
             x"F6",
             x"E6",
             x"F6",
             x"D0",
             x"02",
             x"E6",
             x"F7",
             x"AD",
             x"FD",
             x"FE",
             x"91",
             x"F6",
             x"E6",
             x"F6",
             x"D0",
             x"02",
             x"E6",
             x"F7",
             x"68",
             x"A8",
             x"68",
             x"40",
             x"0F",
             x"23",
             x"F6",
             x"F6",
             x"F6",
             x"F6",
             x"E4",
             x"06",
             x"FE",
             x"FE",
             x"00",
             x"00",
             x"00",
             x"00",
             x"FD",
             x"FE",
             x"0D",
             x"1E",
             x"2F",
             x"4E",
             x"C0",
             x"C0",
             x"C0",
             x"C0",
             x"FE",
             x"FE",
             x"FE",
             x"FE",
             x"FE",
             x"FE",
             x"FE",
             x"FE",
             x"2C",
             x"F8",
             x"FE",
             x"30",
             x"0F",
             x"2C",
             x"FE",
             x"FE",
             x"10",
             x"F6",
             x"A5",
             x"FC",
             x"08",
             x"58",
             x"28",
             x"85",
             x"FC",
             x"4C",
             x"8D",
             x"FE",
             x"AD",
             x"F9",
             x"FE",
             x"60",
             x"68",
             x"85",
             x"FA",
             x"68",
             x"85",
             x"FB",
             x"A0",
             x"00",
             x"E6",
             x"FA",
             x"D0",
             x"02",
             x"E6",
             x"FB",
             x"B1",
             x"FA",
             x"30",
             x"06",
             x"20",
             x"EE",
             x"FF",
             x"4C",
             x"AD",
             x"FE",
             x"6C",
             x"FA",
             x"00",
             x"8D",
             x"FD",
             x"FE",
             x"40",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"00",
             x"00",
             x"00",
             x"00",
             x"00",
             x"00",
             x"00",
             x"00",
             x"00",
             x"00",
             x"00",
             x"00",
             x"00",
             x"00",
             x"00",
             x"00",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"FF",
             x"C4",
             x"FC",
             x"50",
             x"F9",
             x"FD",
             x"FC",
             x"C4",
             x"FC",
             x"D5",
             x"F9",
             x"80",
             x"FA",
             x"0C",
             x"FB",
             x"6D",
             x"F9",
             x"77",
             x"F9",
             x"60",
             x"FC",
             x"D9",
             x"FB",
             x"37",
             x"FC",
             x"43",
             x"FC",
             x"9B",
             x"FC",
             x"19",
             x"FC",
             x"C4",
             x"FC",
             x"88",
             x"F9",
             x"C4",
             x"FC",
             x"C4",
             x"FC",
             x"C4",
             x"FC",
             x"C4",
             x"FC",
             x"C4",
             x"FC",
             x"C4",
             x"FC",
             x"C4",
             x"FC",
             x"88",
             x"F9",
             x"88",
             x"F9",
             x"88",
             x"F9",
             x"36",
             x"80",
             x"FF",
             x"4C",
             x"C4",
             x"FC",
             x"4C",
             x"C4",
             x"FC",
             x"4C",
             x"C4",
             x"FC",
             x"4C",
             x"C4",
             x"FC",
             x"4C",
             x"C4",
             x"FC",
             x"4C",
             x"77",
             x"F9",
             x"4C",
             x"6D",
             x"F9",
             x"6C",
             x"1C",
             x"02",
             x"6C",
             x"1A",
             x"02",
             x"6C",
             x"18",
             x"02",
             x"6C",
             x"16",
             x"02",
             x"6C",
             x"14",
             x"02",
             x"6C",
             x"12",
             x"02",
             x"6C",
             x"10",
             x"02",
             x"C9",
             x"0D",
             x"D0",
             x"07",
             x"A9",
             x"0A",
             x"20",
             x"EE",
             x"FF",
             x"A9",
             x"0D",
             x"6C",
             x"0E",
             x"02",
             x"6C",
             x"0C",
             x"02",
             x"6C",
             x"0A",
             x"02",
             x"6C",
             x"08",
             x"02",
             x"0D",
             x"FE",
             x"00",
             x"F8",
             x"F2",
             x"FC"
    );

begin

    p_rom_bram : process(CLK)
    begin
        if rising_edge(CLK) then
            DATA <= rom(to_integer(unsigned(ADDR)));
        end if;
    end process;

end RTL;
